module adc_sel (
    channel
);

output [4:0] channel;

assign channel = 8;

endmodule
